module button
(
    input wire PIN_2,
    output wire LED
);

assign LED = PIN_2;

endmodule
