module simple;
endmodule

